.title KiCad schematic
P1 NC_01 NC_02 NC_03 +3V3 IN+ GND GND NC_04 Power
P2 NC_05 NC_06 NC_07 NC_08 /A4_SDA_ /A5_SCL_ Analog
P5 NC_09 CONN_01X01
P6 NC_10 CONN_01X01
P7 NC_11 CONN_01X01
P8 NC_12 CONN_01X01
P4 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 Digital
P3 /A5_SCL_ /A4_SDA_ NC_21 GND NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 Digital
U1 Net-_Q1-Pad1_ Net-_Q1-Pad1_ Trigger GND Trigger Net-_Q2-Pad1_ Net-_Q2-Pad1_ IN+ LMV358
R1 GND Trigger 10k
R2 IN+ Net-_D1-Pad2_ 2
R3 IN+ Net-_D1-Pad2_ 2
R4 IN+ Net-_D1-Pad2_ 2
R5 IN+ Net-_D1-Pad2_ 2
C1 IN+ GND 470n
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ LED
Q1 Net-_Q1-Pad1_ GND Net-_D1-Pad1_ DMN3051L
R6 GND Net-_Q1-Pad1_ 10k
C2 IN+ GND 500u
R7 IN+ Net-_D2-Pad2_ 2
R8 IN+ Net-_D2-Pad2_ 2
R9 IN+ Net-_D2-Pad2_ 2
R10 IN+ Net-_D2-Pad2_ 2
D2 Net-_D2-Pad1_ Net-_D2-Pad2_ LED
Q2 Net-_Q2-Pad1_ GND Net-_D2-Pad1_ DMN3051L
C3 IN+ GND 500u
R11 GND Net-_Q2-Pad1_ 10k
.end
